/*
Edited by John lee and Elizabeth Thompson
*/
module hexdriver (input [3:0] val, output logic [6:0] HEX);

	always_comb begin
		case (val)
			4'b0000: HEX = 7'b100_0000; // 0
			4'b0001: HEX = 7'b111_1001; // 1
			4'b0010: HEX = 7'b010_0100; // 2
			4'b0011: HEX = 7'b011_0000; // 3
			4'b0100: HEX = 7'b001_1001; // 4
			
			4'b0101: HEX = 7'b001_0010; // 5 
			
			4'b0110: HEX = 7'b000_0010; // 6
			
			4'b0111: HEX = 7'b111_1000; // 7
			
			4'b1000: HEX = 7'b000_0000; // 8
			
			4'b1001: HEX = 7'b001_1000; // 9 
			4'b1010: HEX = 7'b000_1000; // A 
			
			4'b1011: HEX = 7'b000_0011; // b
			4'b1100: HEX = 7'b100_0110; // C
			4'b1101: HEX = 7'b010_0001; // d
			4'b1110: HEX = 7'b000_0110; // E
			4'b1111: HEX = 7'b000_1110; // F 
			
			//default: HEX = 7'b000_0000;
		endcase
	end
	
	/* your code here */
endmodule
